module ComboDistributor(
  input        clock,
  input        reset,
  output       in_ready, // @[src/main/scala/exercise2/Distributor.scala 27:14]
  input        in_valid, // @[src/main/scala/exercise2/Distributor.scala 27:14]
  input  [7:0] in_bits, // @[src/main/scala/exercise2/Distributor.scala 27:14]
  input  [3:0] dest, // @[src/main/scala/exercise2/Distributor.scala 28:16]
  input        out_0_ready, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output       out_0_valid, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output [7:0] out_0_bits, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  input        out_1_ready, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output       out_1_valid, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output [7:0] out_1_bits, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  input        out_2_ready, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output       out_2_valid, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output [7:0] out_2_bits, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  input        out_3_ready, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output       out_3_valid, // @[src/main/scala/exercise2/Distributor.scala 43:15]
  output [7:0] out_3_bits // @[src/main/scala/exercise2/Distributor.scala 43:15]
);
  wire  _GEN_7 = dest[1] & out_1_ready; // @[src/main/scala/exercise2/Distributor.scala 149:11 140:20]
  wire  allreadyVec_1 = in_valid & _GEN_7; // @[src/main/scala/exercise2/Distributor.scala 140:20 145:4]
  wire  _GEN_3 = dest[0] & out_0_ready; // @[src/main/scala/exercise2/Distributor.scala 149:11 140:20]
  wire  allreadyVec_0 = in_valid & _GEN_3; // @[src/main/scala/exercise2/Distributor.scala 140:20 145:4]
  wire  _GEN_15 = dest[3] & out_3_ready; // @[src/main/scala/exercise2/Distributor.scala 149:11 140:20]
  wire  allreadyVec_3 = in_valid & _GEN_15; // @[src/main/scala/exercise2/Distributor.scala 140:20 145:4]
  wire  _GEN_11 = dest[2] & out_2_ready; // @[src/main/scala/exercise2/Distributor.scala 149:11 140:20]
  wire  allreadyVec_2 = in_valid & _GEN_11; // @[src/main/scala/exercise2/Distributor.scala 140:20 145:4]
  wire [3:0] allready = {allreadyVec_3,allreadyVec_2,allreadyVec_1,allreadyVec_0}; // @[src/main/scala/exercise2/Distributor.scala 134:30]
  wire [7:0] _GEN_2 = dest[0] ? in_bits : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 149:11 139:17 151:25]
  wire [7:0] _GEN_6 = dest[1] ? in_bits : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 149:11 139:17 151:25]
  wire [7:0] _GEN_10 = dest[2] ? in_bits : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 149:11 139:17 151:25]
  wire [7:0] _GEN_14 = dest[3] ? in_bits : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 149:11 139:17 151:25]
  wire  _T_4 = allready == dest; // @[src/main/scala/exercise2/Distributor.scala 158:23]
  assign in_ready = in_valid & _T_4; // @[src/main/scala/exercise2/Distributor.scala 142:12 145:4]
  assign out_0_valid = in_valid & dest[0]; // @[src/main/scala/exercise2/Distributor.scala 138:18 145:4]
  assign out_0_bits = in_valid ? _GEN_2 : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 139:17 145:4]
  assign out_1_valid = in_valid & dest[1]; // @[src/main/scala/exercise2/Distributor.scala 138:18 145:4]
  assign out_1_bits = in_valid ? _GEN_6 : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 139:17 145:4]
  assign out_2_valid = in_valid & dest[2]; // @[src/main/scala/exercise2/Distributor.scala 138:18 145:4]
  assign out_2_bits = in_valid ? _GEN_10 : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 139:17 145:4]
  assign out_3_valid = in_valid & dest[3]; // @[src/main/scala/exercise2/Distributor.scala 138:18 145:4]
  assign out_3_bits = in_valid ? _GEN_14 : 8'h0; // @[src/main/scala/exercise2/Distributor.scala 139:17 145:4]
endmodule
